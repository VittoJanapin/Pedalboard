module distortion (
    CLOCK_50,
    enable,
    left_channel_audio_in,
    right_channel_audio_in,
    left_channel_audio_out,
    right_channel_audio_out,
);

/****************************************************************

                        PORTS                                   
    
*****************************************************************/

input CLOCK_50, enable;
input [31:0] left_channel_audio_in, right_channel_audio_in;
output [31:0] left_channel_audio_out, left_channel_audio_out;

/****************************************************************

                    COMBINATIONAL CIRCUITS                      
    
*****************************************************************/
localparam threshold = 31'b1111111111111;
//lut generated by chatgpt which maps values from 111_111_111_111_111_111 to d5210112

reg [15:0] LUT [0:255] = '{

};
wire [7:0] left_LUT_index;
assign left_LUT_index = left_channel_audio_in[30:23];
wire [7:0] right_LUT_index;
assign right_LUT_index = right_channel_audio_in[30:23];
always @ (*) 
    begin   
        if(~enable) 
        begin
            left_channel_audio_out = left_channel_audio_in;
            right_channel_audio_out = right_channel_audio_in;
        end

        else
        begin
            /***** APPLY DISTORTION LOGIC ******/
            //evaluate the amplitude at different thresholds
            //use lut for with the top 8 bits as index, 
        
            left_channel_audio_out = {left_channel_audio_in[31], LUT[left_LUT_index], 15'b111111111111111};
            right_channel_audio_out = {right_channel_audio_in[31], LUT[left_LUT_INDEX], 15'b111111111111111}
        end
    end

//easy!

